//------------------------------------------------------------------------------------------------------------------------------------------------------------
// WIECLAW Manon
// TP2 IA
// 31.03.2023
//Script permettant de tester l'addition de deux nombres de 16 bits.
//------------------------------------------------------------------------------------------------------------------------------------------------------------



`timescale 1ns / 1ps
module stimulus;
	// Inputs
	reg [15:0] e1 = 16'b0000000000000000;
	reg [15:0] e2 = 16'b0000000000000000;
    reg r0;
   
	// Outputs
	wire [15:0] s;
    wire r1;
	// Instantiate the Unit Under Test (UUT)
	operation16 uut (
		e1 [15:0], 
		e2 [15:0], 
        r0,
		s [15:0],
        r1
	);
 
	initial begin
	$dumpfile("add16bit.vcd");
    $dumpvars(0,stimulus);
		// Initialize Inputs
		e1 = 16'b0000000000000000;
		e2 = 16'b0000000000000000;
        r0 = 0;
 
		#5;

		e1 = 16'b0110000010000001;
		e2 = 16'b0100000100000110;
        r0 = 1;

		#10;

		e1 = 16'b1000001000010011;
		e2 = 16'b0001000010000000;
        r0 = 1;

		#10;

		e1 = 16'b1000100100001000;
		e2 = 16'b1101001101001000;
        r0 = 0;

		#10;
		e1 = 16'b0000000000000000;
		e2 = 16'b0000000000000000;
        r0 = 0;
 
	end  
 
	initial begin
		 $monitor("t=%3d e1=%d, e2=%d, r0=%d, s=%d, r1=%d \n",$time,e1,e2, r0,s,r1);
	end
 
endmodule
 

 
