//------------------------------------------------------------------------------------------------------------------------------------------------------------
// WIECLAW Manon
// TP2 IA
// 31.03.2023
//Script permettant d'effectuer l'addition de deux nombres de 16 bits.
//------------------------------------------------------------------------------------------------------------------------------------------------------------



module operation16(e1, e2, r0, s, r1);

    input [15:0] e1;
    input [15:0] e2;
    input r0; 
    output [15:0] s;
    output r1;
    
   assign  {r1 ,s} = e1 + e2 + r0;
   
endmodule
