//------------------------------------------------------------------------------------------------------------------------------------------------------------
// WIECLAW Manon
// TP2 IA
// 31.03.2023
//Script permettant d'effectuer la multiplication de deux nombres de 16 bits.
//------------------------------------------------------------------------------------------------------------------------------------------------------------


module multiplication16(e1, e2, s);

    input [15:0] e1;
    input [15:0] e2;
     
    output [31:0] s;
    
  
   assign  s = e1 * e2 ;
   
  
endmodule
